interface soc_probe_if(
        input clk, rst
    );

    logic[`RegBus] x3;
    logic[`RegBus] x26;
    logic[`RegBus] x27;

endinterface: soc_probe_if