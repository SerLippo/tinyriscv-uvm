class tinyriscv_config extends uvm_object;

    `uvm_object_utils(tinyriscv_config)

    function new(string name="tinyriscv_config");
        super.new(name);
    endfunction: new

endclass: tinyriscv_config